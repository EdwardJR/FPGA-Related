----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:35:05 07/17/2020 
-- Design Name: 
-- Module Name:    CHAR_TO_DECIMAL - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity CHAR_TO_DECIMAL is
	port(
		CLK 	: in std_logic;
		CHAR	: in std_logic_vector(7 downto 0);
	
	);


end CHAR_TO_DECIMAL;

architecture Behavioral of CHAR_TO_DECIMAL is

begin


end Behavioral;

